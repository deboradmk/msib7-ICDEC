magic
tech sky130A
magscale 1 2
timestamp 1729246295
<< dnwell >>
rect -186 -1162 868 1480
<< nwell >>
rect -186 -1295 868 1613
<< nsubdiff >>
rect -150 1543 -90 1577
rect 772 1543 832 1577
rect -150 1517 -116 1543
rect 798 1517 832 1543
rect -150 -1225 -116 -1199
rect 798 -1225 832 -1199
rect -150 -1259 -90 -1225
rect 772 -1259 832 -1225
<< nsubdiffcont >>
rect -90 1543 772 1577
rect -150 -1199 -116 1517
rect 798 -1199 832 1517
rect -90 -1259 772 -1225
<< poly >>
rect 647 1505 739 1520
rect -19 1488 73 1503
rect -19 1454 -3 1488
rect 31 1454 73 1488
rect -19 1438 73 1454
rect 43 1404 73 1438
rect 647 1471 689 1505
rect 723 1471 739 1505
rect 647 1455 739 1471
rect 647 1404 677 1455
rect -17 792 75 807
rect 133 804 331 909
rect -17 758 -1 792
rect 33 758 75 792
rect -17 742 75 758
rect 45 708 75 742
rect 649 792 741 807
rect 649 758 691 792
rect 725 758 741 792
rect 649 742 741 758
rect 649 708 679 742
rect 134 111 591 213
rect 46 -420 76 -386
rect -16 -436 76 -420
rect -16 -470 0 -436
rect 34 -470 76 -436
rect -16 -485 76 -470
rect 650 -420 680 -386
rect 650 -436 742 -420
rect 650 -470 692 -436
rect 726 -470 742 -436
rect 391 -584 592 -482
rect 650 -485 742 -470
rect 46 -1115 76 -1084
rect -16 -1131 76 -1115
rect -16 -1165 0 -1131
rect 34 -1165 76 -1131
rect -16 -1180 76 -1165
rect 650 -1114 680 -1080
rect 650 -1130 742 -1114
rect 650 -1164 692 -1130
rect 726 -1164 742 -1130
rect 650 -1179 742 -1164
<< polycont >>
rect -3 1454 31 1488
rect 689 1471 723 1505
rect -1 758 33 792
rect 691 758 725 792
rect 0 -470 34 -436
rect 692 -470 726 -436
rect 0 -1165 34 -1131
rect 692 -1164 726 -1130
<< locali >>
rect -150 1543 -90 1577
rect 772 1543 832 1577
rect -150 1517 -116 1543
rect 798 1517 832 1543
rect -19 1454 -3 1488
rect 31 1454 47 1488
rect 673 1471 689 1505
rect 723 1471 739 1505
rect -4 1403 31 1454
rect -3 1400 31 1403
rect 689 1388 724 1471
rect -17 758 -1 792
rect 33 758 49 792
rect 675 758 691 792
rect 725 758 741 792
rect -2 711 33 758
rect -1 708 33 711
rect 691 711 726 758
rect 691 708 725 711
rect 0 -389 34 -386
rect -1 -436 34 -389
rect 692 -389 726 -386
rect 692 -436 727 -389
rect -16 -470 0 -436
rect 34 -470 50 -436
rect 676 -470 692 -436
rect 726 -470 742 -436
rect 0 -1084 34 -1068
rect -1 -1131 34 -1084
rect 692 -1083 726 -1080
rect 692 -1130 727 -1083
rect -16 -1165 0 -1131
rect 34 -1165 50 -1131
rect 676 -1164 692 -1130
rect 726 -1164 742 -1130
rect -150 -1225 -116 -1199
rect 798 -1225 832 -1199
rect -150 -1259 -90 -1225
rect 772 -1259 832 -1225
<< viali >>
rect 689 1543 723 1577
rect -3 1454 31 1488
rect 689 1471 723 1505
rect -1 758 33 792
rect 691 758 725 792
rect 0 -470 34 -436
rect 692 -470 726 -436
rect 0 -1165 34 -1131
rect 692 -1164 726 -1130
rect 0 -1259 34 -1225
<< metal1 >>
rect 677 1577 735 1583
rect 677 1543 689 1577
rect 723 1543 735 1577
rect 678 1505 735 1543
rect -15 1488 43 1494
rect -15 1454 -3 1488
rect 31 1454 43 1488
rect 677 1471 689 1505
rect 723 1471 735 1505
rect 677 1465 735 1471
rect -15 1448 43 1454
rect -10 1403 37 1448
rect -14 1393 130 1403
rect -22 1016 -12 1393
rect 40 1016 130 1393
rect -14 1002 130 1016
rect 340 962 383 1404
rect 683 1400 730 1465
rect 684 1392 726 1400
rect 601 1380 726 1392
rect 601 1016 723 1380
rect 596 962 641 1010
rect 340 914 641 962
rect -13 792 45 798
rect -13 758 -1 792
rect 33 758 45 792
rect -13 752 45 758
rect -8 708 39 752
rect -6 706 41 708
rect -6 700 129 706
rect -7 695 129 700
rect -7 319 79 695
rect 131 319 141 695
rect -7 306 129 319
rect 88 101 175 106
rect 88 95 190 101
rect 87 55 190 95
rect 87 14 122 55
rect -6 -386 130 14
rect -7 -387 99 -386
rect -7 -430 40 -387
rect -12 -436 46 -430
rect -12 -470 0 -436
rect 34 -470 46 -436
rect -12 -476 46 -470
rect 340 -593 383 914
rect 679 792 737 798
rect 679 758 691 792
rect 725 758 737 792
rect 679 752 737 758
rect 685 708 732 752
rect 596 308 732 708
rect 603 267 638 308
rect 556 227 638 267
rect 597 2 733 14
rect 584 -374 594 2
rect 646 -374 733 2
rect 597 -386 733 -374
rect 686 -430 733 -386
rect 680 -436 738 -430
rect 680 -470 692 -436
rect 726 -470 738 -436
rect 680 -476 738 -470
rect 82 -598 383 -593
rect 82 -642 384 -598
rect 82 -683 128 -642
rect 0 -1068 122 -692
rect 340 -1080 383 -642
rect 598 -691 734 -681
rect 598 -1068 683 -691
rect 735 -1068 745 -691
rect 598 -1080 734 -1068
rect -7 -1125 40 -1080
rect 598 -1081 733 -1080
rect 686 -1124 733 -1081
rect -12 -1131 46 -1125
rect -12 -1165 0 -1131
rect 34 -1165 46 -1131
rect -12 -1225 46 -1165
rect 680 -1130 738 -1124
rect 680 -1164 692 -1130
rect 726 -1164 738 -1130
rect 680 -1170 738 -1164
rect -12 -1259 0 -1225
rect 34 -1259 46 -1225
rect -12 -1265 46 -1259
<< via1 >>
rect -12 1016 40 1393
rect 79 319 131 695
rect 594 -374 646 2
rect 683 -1068 735 -691
<< metal2 >>
rect -8 1403 40 1489
rect -12 1393 40 1403
rect -12 1006 40 1016
rect -8 900 40 1006
rect -12 891 44 900
rect 685 893 733 894
rect -12 826 44 835
rect 669 833 678 893
rect 738 833 747 893
rect -8 -487 40 826
rect 79 695 131 705
rect 79 309 131 319
rect 85 180 120 309
rect 85 153 638 180
rect 86 146 638 153
rect 604 12 638 146
rect 594 2 646 12
rect 594 -384 646 -374
rect -15 -492 47 -487
rect 685 -488 733 833
rect -25 -495 55 -492
rect -25 -555 -14 -495
rect 46 -555 55 -495
rect -25 -557 55 -555
rect 685 -497 741 -488
rect -15 -566 47 -557
rect 685 -562 741 -553
rect 687 -681 732 -562
rect 683 -691 735 -681
rect 683 -1078 735 -1068
rect 687 -1080 732 -1078
<< via2 >>
rect -12 835 44 891
rect 678 833 738 893
rect -14 -555 46 -495
rect 685 -553 741 -497
<< metal3 >>
rect -17 893 49 896
rect 673 893 743 898
rect -17 891 678 893
rect -17 835 -12 891
rect 44 835 678 891
rect -17 833 678 835
rect 738 833 743 893
rect -17 830 49 833
rect 673 828 743 833
rect -19 -495 51 -490
rect 680 -495 746 -492
rect -19 -555 -14 -495
rect 46 -497 746 -495
rect 46 -553 685 -497
rect 741 -553 746 -497
rect 46 -555 746 -553
rect -19 -560 51 -555
rect 680 -558 746 -555
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729134042
transform 1 0 665 0 1 -880
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729134042
transform 1 0 60 0 1 508
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729134042
transform 1 0 61 0 1 -880
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_3
timestamp 1729134042
transform 1 0 61 0 1 -186
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729134042
transform 1 0 665 0 1 -186
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729134042
transform 1 0 664 0 1 508
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729134042
transform 1 0 662 0 1 1204
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729134042
transform 1 0 58 0 1 1204
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729147639
transform 1 0 360 0 1 1204
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729147639
transform 1 0 362 0 1 508
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729147639
transform 1 0 363 0 1 -186
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729147639
transform 1 0 363 0 1 -880
box -323 -300 323 300
<< labels >>
flabel metal1 616 248 616 248 0 FreeSans 480 0 0 0 D2
port 8 nsew
flabel metal2 101 159 101 159 0 FreeSans 480 0 0 0 D1
port 10 nsew
flabel metal2 708 102 708 102 0 FreeSans 480 0 0 0 D5
port 12 nsew
flabel metal1 709 1528 709 1528 0 FreeSans 480 0 0 0 VDD
port 14 nsew
<< end >>
