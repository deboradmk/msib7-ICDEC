magic
tech sky130A
magscale 1 2
timestamp 1729408806
<< nwell >>
rect -176 -305 622 2014
<< pmos >>
rect 410 1408 440 1410
rect 410 972 440 974
<< pdiff >>
rect 401 1408 410 1410
rect 440 1408 498 1410
rect 404 972 410 974
rect 440 972 498 974
<< nsubdiff >>
rect -140 1944 -80 1978
rect 526 1944 586 1978
rect -140 1701 -106 1944
rect 552 1701 586 1944
rect -140 -235 -106 7
rect 552 -235 586 7
rect -140 -269 -80 -235
rect 526 -269 586 -235
<< nsubdiffcont >>
rect -80 1944 526 1978
rect -140 7 -106 1701
rect 552 7 586 1701
rect -80 -269 526 -235
<< poly >>
rect 6 1377 36 1408
rect -56 1361 36 1377
rect -56 1327 -40 1361
rect -6 1327 36 1361
rect -56 1311 36 1327
rect 410 1377 440 1408
rect 410 1361 502 1377
rect 410 1327 452 1361
rect 486 1327 502 1361
rect 410 1311 502 1327
rect 6 941 36 970
rect -56 925 36 941
rect -56 891 -40 925
rect -6 891 36 925
rect 410 941 440 972
rect 410 925 502 941
rect -56 875 36 891
rect -56 817 36 833
rect 94 817 194 891
rect 253 818 353 892
rect 410 891 452 925
rect 486 891 502 925
rect 410 875 502 891
rect 410 817 502 833
rect -56 783 -40 817
rect -6 783 36 817
rect -56 767 36 783
rect 6 736 36 767
rect 410 783 452 817
rect 486 783 502 817
rect 410 767 502 783
rect 410 736 440 767
rect -56 382 36 398
rect -56 348 -40 382
rect -6 348 36 382
rect -56 332 36 348
rect 6 279 36 332
rect 410 381 502 397
rect 410 347 452 381
rect 486 347 502 381
rect 410 331 502 347
rect 410 279 440 331
<< polycont >>
rect -40 1327 -6 1361
rect 452 1327 486 1361
rect -40 891 -6 925
rect 452 891 486 925
rect -40 783 -6 817
rect 452 783 486 817
rect -40 348 -6 382
rect 452 347 486 381
<< locali >>
rect -140 1944 -80 1978
rect 526 1944 586 1978
rect -140 1701 -106 1944
rect 552 1701 586 1944
rect 452 1569 486 1610
rect -40 1406 -6 1408
rect -41 1361 -6 1406
rect 48 1404 49 1408
rect 452 1406 486 1410
rect 452 1361 487 1406
rect -56 1327 -40 1361
rect -6 1327 10 1361
rect 436 1327 452 1361
rect 486 1327 502 1361
rect 452 1134 486 1170
rect -40 970 -6 997
rect -41 925 -6 970
rect 48 969 54 971
rect 452 970 486 974
rect 452 925 487 970
rect -56 891 -40 925
rect -6 891 10 925
rect 436 891 452 925
rect 486 891 502 925
rect -56 783 -40 817
rect -6 783 10 817
rect 436 783 452 817
rect 486 783 502 817
rect -41 700 -6 783
rect 452 736 486 783
rect -56 348 -40 382
rect -6 348 10 382
rect -40 277 -6 348
rect 436 347 452 381
rect 486 347 502 381
rect 452 256 486 347
rect -140 -235 -106 7
rect 552 -235 586 7
rect -140 -269 -80 -235
rect 526 -269 586 -235
<< viali >>
rect 106 1978 248 1979
rect 106 1944 248 1978
rect -40 1327 -6 1361
rect 452 1327 486 1361
rect -40 891 -6 925
rect 452 891 486 925
rect -40 783 -6 817
rect 452 783 486 817
rect -40 348 -6 382
rect 452 347 486 381
<< metal1 >>
rect 94 1979 260 1985
rect 94 1944 106 1979
rect 248 1944 260 1979
rect 94 1938 260 1944
rect 471 1914 523 1920
rect -5 1865 471 1910
rect -5 1607 47 1865
rect 471 1856 523 1862
rect 487 1779 493 1790
rect 129 1750 493 1779
rect 129 1657 158 1750
rect 487 1738 493 1750
rect 545 1738 551 1790
rect -45 1586 82 1607
rect -46 1426 82 1586
rect 390 1584 400 1610
rect 187 1483 197 1535
rect 249 1483 259 1535
rect -45 1408 82 1426
rect 366 1424 400 1584
rect 390 1409 400 1424
rect 452 1563 493 1610
rect 452 1424 492 1563
rect 452 1410 462 1424
rect 452 1409 493 1410
rect 401 1408 404 1409
rect -47 1407 82 1408
rect -47 1367 0 1407
rect -52 1361 6 1367
rect -52 1327 -40 1361
rect -6 1327 6 1361
rect -52 1321 6 1327
rect 270 1318 280 1370
rect 332 1318 342 1370
rect 446 1367 493 1409
rect 440 1361 498 1367
rect 440 1327 452 1361
rect 486 1327 498 1361
rect 440 1321 498 1327
rect 492 1262 544 1268
rect 102 1208 112 1260
rect 164 1208 174 1260
rect 302 1219 492 1253
rect 492 1204 544 1210
rect -62 970 -52 1171
rect 0 1164 10 1171
rect 0 1004 84 1164
rect 453 1159 463 1161
rect 445 1152 463 1159
rect 185 1042 195 1102
rect 255 1042 265 1102
rect 370 1064 463 1152
rect 0 970 10 1004
rect 362 984 463 1064
rect 522 984 532 1161
rect 362 976 500 984
rect -47 931 0 970
rect -52 925 6 931
rect -52 891 -40 925
rect -6 891 6 925
rect -52 885 6 891
rect 440 925 500 976
rect 440 891 452 925
rect 486 910 500 925
rect 486 891 498 910
rect 440 885 498 891
rect -52 817 6 823
rect -52 783 -40 817
rect -6 783 6 817
rect -52 777 6 783
rect 440 817 498 823
rect 440 783 452 817
rect 486 783 498 817
rect 440 777 498 783
rect -47 738 0 777
rect -62 537 -52 738
rect 0 732 10 738
rect 445 736 491 777
rect 0 538 80 732
rect 455 723 465 725
rect 450 704 465 723
rect 185 605 195 665
rect 255 605 265 665
rect 360 548 465 704
rect 524 548 534 725
rect 360 544 486 548
rect 0 537 10 538
rect 494 498 546 504
rect 100 446 110 498
rect 162 446 172 498
rect 303 455 494 489
rect 494 440 546 446
rect -52 382 6 388
rect -52 348 -40 382
rect -6 348 6 382
rect 118 367 194 381
rect -52 342 6 348
rect 169 347 194 367
rect -47 301 -1 342
rect 273 338 283 390
rect 335 338 345 390
rect 440 381 498 387
rect 440 347 452 381
rect 486 347 498 381
rect 440 341 498 347
rect 445 301 491 341
rect -47 264 47 301
rect 389 272 399 301
rect -47 259 78 264
rect -30 104 78 259
rect 185 169 195 229
rect 255 169 265 229
rect 368 112 399 272
rect -5 -155 47 104
rect 389 100 399 112
rect 451 272 491 301
rect 451 112 494 272
rect 451 100 461 112
rect 130 -32 160 53
rect 494 -21 546 -15
rect 130 -62 494 -32
rect 494 -79 546 -73
rect 467 -147 527 -141
rect 384 -155 467 -154
rect -5 -200 467 -155
rect -5 -201 47 -200
rect 467 -213 527 -207
<< via1 >>
rect 471 1862 523 1914
rect 493 1738 545 1790
rect 197 1483 249 1535
rect 400 1409 452 1610
rect 280 1318 332 1370
rect 112 1208 164 1260
rect 492 1210 544 1262
rect -52 970 0 1171
rect 195 1042 255 1102
rect 463 984 522 1161
rect -52 537 0 738
rect 195 605 255 665
rect 465 548 524 725
rect 110 446 162 498
rect 494 446 546 498
rect 283 338 335 390
rect 195 169 255 229
rect 399 100 451 301
rect 494 -73 546 -21
rect 467 -207 527 -147
<< metal2 >>
rect 467 1918 527 1927
rect 465 1862 467 1914
rect 527 1862 529 1914
rect 467 1849 527 1858
rect -51 1759 448 1799
rect -51 1702 -6 1759
rect -51 1181 -5 1702
rect 403 1620 448 1759
rect 493 1790 545 1796
rect 493 1732 545 1738
rect 400 1610 452 1620
rect 195 1537 251 1547
rect 195 1471 251 1481
rect 400 1399 452 1409
rect 280 1370 332 1380
rect 280 1311 332 1318
rect 120 1308 332 1311
rect 120 1275 323 1308
rect 120 1270 164 1275
rect 112 1260 164 1270
rect 504 1262 533 1732
rect 486 1210 492 1262
rect 544 1210 550 1262
rect 112 1198 164 1208
rect -52 1171 0 1181
rect 463 1161 522 1171
rect 195 1102 255 1112
rect 195 1032 255 1042
rect 463 974 522 984
rect -52 960 0 970
rect -51 748 -5 960
rect -52 738 0 748
rect 465 725 524 735
rect 195 665 255 675
rect 195 595 255 605
rect 465 538 524 548
rect -52 527 0 537
rect -51 -43 -5 527
rect 110 498 162 508
rect 488 446 494 498
rect 546 446 552 498
rect 110 445 162 446
rect 110 436 330 445
rect 115 404 330 436
rect 283 400 330 404
rect 283 390 335 400
rect 283 328 335 338
rect 399 301 451 311
rect 195 229 255 239
rect 195 159 255 169
rect 399 90 451 100
rect 401 -43 446 90
rect 505 -21 535 446
rect -51 -81 447 -43
rect 488 -73 494 -21
rect 546 -73 552 -21
rect 469 -147 525 -140
rect 461 -207 467 -147
rect 527 -207 533 -147
rect 469 -214 525 -207
<< via2 >>
rect 467 1914 527 1918
rect 467 1862 471 1914
rect 471 1862 523 1914
rect 523 1862 527 1914
rect 467 1858 527 1862
rect 195 1535 251 1537
rect 195 1483 197 1535
rect 197 1483 249 1535
rect 249 1483 251 1535
rect 195 1481 251 1483
rect 195 1042 255 1102
rect 463 984 522 1161
rect 195 605 255 665
rect 465 548 524 725
rect 195 169 255 229
rect 469 -205 525 -149
<< metal3 >>
rect 462 1918 532 1923
rect 462 1858 467 1918
rect 527 1858 532 1918
rect 462 1853 532 1858
rect 185 1537 261 1542
rect 185 1481 195 1537
rect 251 1481 261 1537
rect 185 1476 261 1481
rect 195 1107 255 1476
rect 467 1166 527 1853
rect 453 1161 532 1166
rect 185 1102 265 1107
rect 185 1042 195 1102
rect 255 1042 265 1102
rect 185 1037 265 1042
rect 195 670 255 1037
rect 453 984 463 1161
rect 522 984 532 1161
rect 453 979 532 984
rect 467 730 527 979
rect 455 725 534 730
rect 185 665 265 670
rect 185 605 195 665
rect 255 605 265 665
rect 185 600 265 605
rect 195 234 255 600
rect 455 548 465 725
rect 524 548 534 725
rect 455 543 534 548
rect 185 229 265 234
rect 185 169 195 229
rect 255 169 265 229
rect 185 164 265 169
rect 467 -144 527 543
rect 464 -149 530 -144
rect 464 -205 469 -149
rect 525 -205 530 -149
rect 464 -210 530 -205
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729355162
transform 1 0 425 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729355162
transform 1 0 21 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729355162
transform 1 0 21 0 1 636
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729355162
transform 1 0 21 0 1 1072
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1729355162
transform 1 0 21 0 1 1508
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1729355162
transform 1 0 425 0 1 1508
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1729355162
transform 1 0 425 0 1 1072
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_7
timestamp 1729355162
transform 1 0 425 0 1 636
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_BHV229  sky130_fd_pr__pfet_01v8_BHV229_0
timestamp 1729355162
transform 1 0 223 0 1 854
box -223 -854 223 854
<< labels >>
flabel viali 198 1958 198 1958 0 FreeSans 800 0 0 0 VDD
port 0 nsew
flabel metal2 -30 1770 -30 1770 0 FreeSans 800 0 0 0 D6
port 4 nsew
flabel metal1 383 1236 383 1236 0 FreeSans 800 0 0 0 VIP
port 12 nsew
flabel metal2 149 418 149 418 0 FreeSans 800 0 0 0 VIN
port 14 nsew
flabel metal1 404 -176 406 -176 0 FreeSans 800 0 0 0 OUT
port 16 nsew
flabel metal3 222 1356 222 1356 0 FreeSans 800 0 0 0 D5
port 18 nsew
<< end >>
