magic
tech sky130A
magscale 1 2
timestamp 1729344768
<< psubdiff >>
rect -290 831 -211 865
rect 1530 831 1590 865
rect -290 805 -256 831
rect 1556 805 1590 831
rect -290 -38 -256 -12
rect 1556 -38 1590 -12
rect -290 -72 -211 -38
rect 1530 -72 1590 -38
<< psubdiffcont >>
rect -211 831 1530 865
rect -290 -12 -256 805
rect 1556 -12 1590 805
rect -211 -72 1530 -38
<< poly >>
rect -161 779 -95 795
rect -161 745 -145 779
rect -111 745 -95 779
rect -161 729 -95 745
rect 1368 779 1434 795
rect 1368 745 1384 779
rect 1418 745 1434 779
rect 1368 729 1434 745
rect 1386 706 1416 729
rect 58 366 1214 428
rect -144 66 -114 106
rect -162 50 -96 66
rect 1386 62 1416 88
rect -162 16 -146 50
rect -112 16 -96 50
rect -162 0 -96 16
rect 1368 46 1434 62
rect 1368 12 1384 46
rect 1418 12 1434 46
rect 1368 -4 1434 12
<< polycont >>
rect -145 745 -111 779
rect 1384 745 1418 779
rect -146 16 -112 50
rect 1384 12 1418 46
<< locali >>
rect -290 831 -211 865
rect 1530 831 1590 865
rect -290 805 -256 831
rect 1556 805 1590 831
rect -194 782 -152 784
rect -104 782 -62 784
rect -194 779 -62 782
rect -194 745 -145 779
rect -111 745 -62 779
rect -194 734 -62 745
rect -194 690 -152 734
rect -104 690 -62 734
rect 1336 779 1466 784
rect 1336 745 1384 779
rect 1418 745 1466 779
rect 1336 736 1466 745
rect 1336 690 1378 736
rect 1424 690 1466 736
rect -194 64 -152 110
rect -106 64 -64 106
rect -194 50 -64 64
rect -194 16 -146 50
rect -112 16 -64 50
rect -106 12 -64 16
rect 1334 54 1376 100
rect 1424 54 1466 102
rect 1334 46 1466 54
rect 1334 12 1384 46
rect 1418 12 1466 46
rect 1334 8 1466 12
rect 1334 6 1438 8
rect -290 -38 -256 -12
rect 1556 -38 1590 -12
rect -290 -72 -211 -38
rect 1530 -72 1590 -38
<< viali >>
rect 595 865 676 870
rect 595 832 676 865
rect -145 745 -111 779
rect 1384 745 1418 779
rect -146 16 -112 50
rect 1384 12 1418 46
rect 591 -38 674 -25
rect 591 -72 674 -38
rect 591 -83 674 -72
<< metal1 >>
rect 583 870 690 876
rect 583 859 595 870
rect 270 832 595 859
rect 676 859 690 870
rect 676 832 1008 859
rect 270 826 1008 832
rect -189 779 -67 785
rect -189 745 -145 779
rect -111 745 -67 779
rect -189 739 -67 745
rect -189 700 -155 739
rect -101 700 -67 739
rect -194 510 52 700
rect 12 474 46 510
rect 12 428 74 474
rect -102 282 -68 292
rect -194 281 52 282
rect -194 229 -112 281
rect -60 229 52 281
rect -194 92 52 229
rect -190 56 -156 92
rect -102 56 -68 92
rect -190 50 -68 56
rect -190 16 -146 50
rect -112 16 -68 50
rect -190 10 -68 16
rect 270 -29 300 826
rect 585 706 690 826
rect 344 474 378 525
rect 344 428 406 474
rect 328 100 338 152
rect 390 100 400 152
rect 579 100 693 706
rect 872 642 882 694
rect 934 642 944 694
rect 865 320 928 366
rect 894 268 928 320
rect 579 -19 685 100
rect 579 -25 686 -19
rect 579 -29 591 -25
rect 270 -62 591 -29
rect 579 -83 591 -62
rect 674 -29 686 -25
rect 977 -28 1008 826
rect 1340 779 1462 785
rect 1340 745 1384 779
rect 1418 745 1462 779
rect 1340 739 1462 745
rect 1340 706 1374 739
rect 1428 706 1462 739
rect 1220 570 1466 700
rect 1220 518 1331 570
rect 1383 518 1466 570
rect 1220 510 1466 518
rect 1340 502 1374 510
rect 1197 320 1260 366
rect 1226 286 1260 320
rect 1224 96 1470 286
rect 1340 52 1374 88
rect 1428 52 1462 88
rect 1340 46 1462 52
rect 1340 12 1384 46
rect 1418 12 1462 46
rect 1340 6 1462 12
rect 969 -29 1008 -28
rect 674 -62 1008 -29
rect 674 -83 686 -62
rect 579 -89 686 -83
<< via1 >>
rect -112 229 -60 281
rect 338 100 390 152
rect 882 642 934 694
rect 1331 518 1383 570
<< metal2 >>
rect 882 694 934 704
rect 339 416 391 417
rect 882 416 934 642
rect 1331 570 1383 580
rect 1331 416 1383 518
rect -112 381 1383 416
rect -112 281 -60 381
rect -112 219 -60 229
rect 339 162 391 381
rect 338 153 391 162
rect 338 152 390 153
rect 338 90 390 100
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1729327062
transform 1 0 1401 0 1 188
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1729327062
transform 1 0 -129 0 1 188
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1729327062
transform 1 0 -128 0 1 606
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1729327062
transform 1 0 1401 0 1 606
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_C77M8X  sky130_fd_pr__nfet_01v8_C77M8X_0
timestamp 1729327062
transform 1 0 636 0 1 397
box -636 -397 636 397
<< labels >>
flabel space 137 611 137 611 0 FreeSans 320 0 0 0 m8
flabel space 471 600 471 602 0 FreeSans 320 0 0 0 m8
flabel space 788 599 788 599 0 FreeSans 320 0 0 0 m9
flabel space 1124 605 1124 605 0 FreeSans 320 0 0 0 m9
flabel space 137 196 137 196 0 FreeSans 320 0 0 0 m9
flabel space 464 184 464 184 0 FreeSans 320 0 0 0 m9
flabel space 802 180 802 180 0 FreeSans 320 0 0 0 m8
flabel space 1136 182 1136 182 0 FreeSans 320 0 0 0 m8
flabel metal1 25 607 25 607 0 FreeSans 320 0 0 0 d8
flabel space 364 607 364 607 0 FreeSans 320 0 0 0 d8
flabel space 577 603 577 603 0 FreeSans 320 0 0 0 s
flabel metal1 690 603 690 603 0 FreeSans 320 0 0 0 s
flabel space 1027 603 1027 603 0 FreeSans 320 0 0 0 s
flabel space 244 605 244 605 0 FreeSans 320 0 0 0 s
flabel metal1 1244 601 1244 601 0 FreeSans 320 0 0 0 d9
flabel metal1 23 188 23 188 0 FreeSans 320 0 0 0 d9
flabel space 915 184 915 184 0 FreeSans 320 0 0 0 d8
flabel space 1025 184 1025 184 0 FreeSans 320 0 0 0 s
flabel space 575 186 575 186 0 FreeSans 320 0 0 0 s
flabel metal1 690 184 690 184 0 FreeSans 320 0 0 0 s
flabel space 248 186 248 186 0 FreeSans 320 0 0 0 s
flabel metal1 1243 187 1243 187 0 FreeSans 320 0 0 0 d8
flabel metal1 1297 210 1297 210 0 FreeSans 1120 0 0 0 d8
port 1 nsew
flabel metal1 1295 609 1295 609 0 FreeSans 1120 0 0 0 d9
port 2 nsew
flabel metal1 638 761 638 761 0 FreeSans 1120 0 0 0 gnd
port 4 nsew
flabel metal2 360 188 360 188 0 FreeSans 320 0 0 0 d9
<< end >>
