magic
tech sky130A
magscale 1 2
timestamp 1729346748
<< psubdiff >>
rect -386 1226 -326 1260
rect 1106 1226 1166 1260
rect -386 1200 -352 1226
rect 1132 1200 1166 1226
rect -386 -38 -352 -12
rect 1132 -38 1166 -12
rect -386 -72 -326 -38
rect 1106 -72 1166 -38
<< psubdiffcont >>
rect -326 1226 1106 1260
rect -386 -12 -352 1200
rect 1132 -12 1166 1200
rect -326 -72 1106 -38
<< poly >>
rect -240 679 -210 705
rect -302 663 -210 679
rect -302 629 -286 663
rect -252 629 -210 663
rect 990 681 1020 707
rect 990 665 1082 681
rect 990 631 1032 665
rect 1066 631 1082 665
rect -302 613 -236 629
rect 57 576 724 619
rect 1016 615 1082 631
rect -239 62 -209 88
rect -301 46 -209 62
rect -301 12 -285 46
rect -251 12 -209 46
rect 989 59 1019 101
rect 989 43 1081 59
rect -301 -4 -235 12
rect 989 9 1031 43
rect 1065 9 1081 43
rect 1015 -7 1081 9
<< polycont >>
rect -286 629 -252 663
rect 1032 631 1066 665
rect -285 12 -251 46
rect 1031 9 1065 43
<< locali >>
rect -386 1226 -326 1260
rect 1106 1226 1166 1260
rect -386 1200 -352 1226
rect 1132 1200 1166 1226
rect -286 663 -252 722
rect 1032 665 1066 723
rect -302 629 -286 663
rect -252 629 -236 663
rect 1016 631 1032 665
rect 1066 631 1082 665
rect 1032 630 1066 631
rect -285 46 -251 104
rect -301 12 -285 46
rect -251 12 -235 46
rect 1031 43 1065 106
rect 1015 9 1031 43
rect 1065 9 1081 43
rect -386 -38 -352 -12
rect 1132 -38 1166 -12
rect -386 -72 -326 -38
rect 1106 -72 1166 -38
<< viali >>
rect 350 1226 384 1260
rect -286 629 -252 663
rect 1032 631 1066 665
rect -285 12 -251 46
rect 1031 9 1065 43
rect 384 -72 418 -38
<< metal1 >>
rect 338 1260 396 1266
rect 338 1226 350 1260
rect 384 1226 396 1260
rect 338 1220 396 1226
rect -292 706 52 1105
rect 350 1097 384 1220
rect 297 1069 384 1097
rect -292 669 -246 706
rect 12 674 46 706
rect 264 705 396 746
rect 459 707 469 1107
rect 523 707 533 1107
rect 730 1103 1074 1106
rect 730 714 802 1103
rect 936 714 1074 1103
rect 730 707 1074 714
rect -298 663 -240 669
rect -298 629 -286 663
rect -252 629 -240 663
rect -298 623 -240 629
rect 12 628 74 674
rect 355 656 396 705
rect 1026 671 1072 707
rect 1020 665 1078 671
rect 328 538 444 656
rect 1020 631 1032 665
rect 1066 631 1078 665
rect 1020 625 1078 631
rect 386 487 423 538
rect 702 521 776 567
rect 730 488 776 521
rect -291 484 53 487
rect -291 95 -148 484
rect -14 375 53 484
rect -13 242 53 375
rect -14 95 53 242
rect -291 88 53 95
rect -291 52 -245 88
rect 252 87 262 487
rect 316 87 326 487
rect 386 450 518 487
rect 384 128 477 131
rect 384 101 512 128
rect -297 46 -239 52
rect -297 12 -285 46
rect -251 12 -239 46
rect -297 6 -239 12
rect 384 -32 418 101
rect 730 89 1074 488
rect 1025 49 1071 89
rect 1019 43 1077 49
rect 1019 9 1031 43
rect 1065 9 1077 43
rect 1019 3 1077 9
rect 372 -38 430 -32
rect 372 -72 384 -38
rect 418 -72 430 -38
rect 372 -78 430 -72
<< via1 >>
rect 469 707 523 1107
rect 802 714 936 1103
rect -148 375 -14 484
rect -148 242 -13 375
rect -148 95 -14 242
rect 262 87 316 487
<< metal2 >>
rect 458 1114 523 1117
rect 458 1107 533 1114
rect 819 1113 923 1120
rect 458 707 469 1107
rect 523 707 533 1107
rect 458 652 533 707
rect 802 1110 936 1113
rect 802 1103 819 1110
rect 923 1103 936 1110
rect 802 710 819 714
rect 923 710 936 714
rect 802 704 936 710
rect 819 700 923 704
rect 255 570 534 652
rect -132 494 -28 497
rect -148 487 -14 494
rect -148 484 -132 487
rect -28 484 -14 487
rect 256 487 326 570
rect -14 375 -13 385
rect -14 232 -13 242
rect -148 87 -132 95
rect -28 87 -14 95
rect -148 85 -14 87
rect 256 87 262 487
rect 316 87 326 487
rect -132 77 -28 85
rect 256 79 326 87
rect 262 77 326 79
<< via2 >>
rect 819 1103 923 1110
rect 819 714 923 1103
rect 819 710 923 714
rect -132 484 -28 487
rect -132 95 -28 484
rect -132 87 -28 95
<< metal3 >>
rect 809 1110 933 1115
rect 809 732 819 1110
rect 808 710 819 732
rect 923 710 933 1110
rect 808 705 933 710
rect 808 653 930 705
rect -133 543 930 653
rect -133 492 -17 543
rect -142 487 -17 492
rect -142 87 -132 487
rect -28 468 -17 487
rect -28 87 -18 468
rect -142 82 -18 87
use sky130_fd_pr__nfet_01v8_4HFSKE  sky130_fd_pr__nfet_01v8_4HFSKE_0
timestamp 1729258563
transform 1 0 -225 0 1 905
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_4HFSKE  sky130_fd_pr__nfet_01v8_4HFSKE_1
timestamp 1729258563
transform 1 0 1005 0 1 907
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_4HFSKE  sky130_fd_pr__nfet_01v8_4HFSKE_2
timestamp 1729258563
transform 1 0 1004 0 1 289
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_4HFSKE  sky130_fd_pr__nfet_01v8_4HFSKE_3
timestamp 1729258563
transform 1 0 -224 0 1 288
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_ZY4669  sky130_fd_pr__nfet_01v8_ZY4669_0
timestamp 1729258563
transform 1 0 624 0 1 598
box -158 -597 158 597
use sky130_fd_pr__nfet_01v8_ZY4669  sky130_fd_pr__nfet_01v8_ZY4669_1
timestamp 1729258563
transform 1 0 158 0 1 597
box -158 -597 158 597
<< labels >>
flabel metal1 364 1173 364 1173 0 FreeSans 800 0 0 0 GND
port 0 nsew
flabel metal1 27 684 27 684 0 FreeSans 800 0 0 0 D3
port 1 nsew
flabel metal3 859 659 859 659 0 FreeSans 800 0 0 0 D4
port 3 nsew
flabel metal2 498 678 498 678 0 FreeSans 800 0 0 0 RS
port 5 nsew
<< end >>
