magic
tech sky130A
magscale 1 2
timestamp 1729337773
use nmoscss  nmoscss_0
timestamp 1729337349
transform 1 0 290 0 1 89
box -290 -89 1590 876
<< labels >>
flabel space 924 30 924 30 0 FreeSans 1600 0 0 0 gnd
port 0 nsew
flabel space 1586 292 1586 292 0 FreeSans 1600 0 0 0 d8
port 1 nsew
flabel space 260 288 260 288 0 FreeSans 1600 0 0 0 d9
port 2 nsew
<< end >>
