magic
tech sky130A
magscale 1 2
timestamp 1729091380
<< viali >>
rect 617 1032 718 1068
rect 1324 1042 1425 1078
rect 2010 1036 2111 1072
rect 613 13 724 47
rect 1323 21 1433 56
rect 2004 16 2114 51
<< metal1 >>
rect 413 1078 2426 1091
rect 413 1068 1324 1078
rect 413 1032 617 1068
rect 718 1042 1324 1068
rect 1425 1072 2426 1078
rect 1425 1042 2010 1072
rect 718 1036 2010 1042
rect 2111 1036 2426 1072
rect 718 1032 2426 1036
rect 413 1022 2426 1032
rect 2278 572 2424 580
rect 385 559 531 567
rect 385 506 404 559
rect 500 552 531 559
rect 500 516 670 552
rect 774 524 1373 559
rect 1482 526 2060 557
rect 2278 556 2304 572
rect 2158 524 2304 556
rect 2278 519 2304 524
rect 2400 519 2424 572
rect 500 506 531 516
rect 2278 508 2424 519
rect 385 495 531 506
rect 395 56 2345 76
rect 395 47 1323 56
rect 395 13 613 47
rect 724 21 1323 47
rect 1433 51 2345 56
rect 1433 21 2004 51
rect 724 16 2004 21
rect 2114 16 2345 51
rect 724 13 2345 16
rect 395 -15 2345 13
<< via1 >>
rect 404 506 500 559
rect 2304 519 2400 572
<< metal2 >>
rect 2279 572 2425 584
rect 2279 568 2304 572
rect 383 559 2304 568
rect 383 506 404 559
rect 500 519 2304 559
rect 2400 519 2425 572
rect 500 510 2425 519
rect 500 506 529 510
rect 2279 509 2425 510
rect 383 493 529 506
use iinverter  iinverter_0 ~/project1
timestamp 1728982223
transform 1 0 513 0 1 -31
box -53 9 369 1135
use iinverter  iinverter_1
timestamp 1728982223
transform 1 0 1217 0 1 -23
box -53 9 369 1135
use iinverter  iinverter_2
timestamp 1728982223
transform 1 0 1901 0 1 -28
box -53 9 369 1135
<< labels >>
flabel metal1 1037 1058 1037 1058 0 FreeSans 320 0 0 0 VVDD
port 0 nsew
flabel metal2 1652 535 1652 535 0 FreeSans 320 0 0 0 OUT
port 1 nsew
flabel metal1 956 22 956 22 0 FreeSans 320 0 0 0 VGND
port 3 nsew
<< end >>
