magic
tech sky130A
magscale 1 2
timestamp 1729337349
<< psubdiff >>
rect -290 831 -211 865
rect 1530 831 1590 865
rect -290 805 -256 831
rect 1556 805 1590 831
rect -290 -38 -256 -12
rect 1556 -38 1590 -12
rect -290 -72 -211 -38
rect 1530 -72 1590 -38
<< psubdiffcont >>
rect -211 831 1530 865
rect -290 -12 -256 805
rect 1556 -12 1590 805
rect -211 -72 1530 -38
<< poly >>
rect -161 779 -95 795
rect -161 745 -145 779
rect -111 745 -95 779
rect -161 729 -95 745
rect 1368 779 1434 795
rect 1368 745 1384 779
rect 1418 745 1434 779
rect 1368 729 1434 745
rect 1386 706 1416 729
rect 58 366 1214 428
rect -144 66 -114 106
rect -162 50 -96 66
rect 1386 62 1416 88
rect -162 16 -146 50
rect -112 16 -96 50
rect -162 0 -96 16
rect 1368 46 1434 62
rect 1368 12 1384 46
rect 1418 12 1434 46
rect 1368 -4 1434 12
<< polycont >>
rect -145 745 -111 779
rect 1384 745 1418 779
rect -146 16 -112 50
rect 1384 12 1418 46
<< locali >>
rect -290 831 -211 865
rect 1530 831 1590 865
rect -290 805 -256 831
rect 1556 805 1590 831
rect -161 745 -145 779
rect -111 745 -95 779
rect 1368 745 1384 779
rect 1418 745 1434 779
rect 1340 706 1374 710
rect 1428 706 1462 710
rect -190 88 -156 92
rect -102 88 -68 92
rect -162 16 -146 50
rect -112 16 -96 50
rect 1368 12 1384 46
rect 1418 12 1434 46
rect -290 -38 -256 -12
rect 1556 -38 1590 -12
rect -290 -72 -211 -38
rect 1530 -72 1590 -38
<< viali >>
rect 595 865 676 870
rect 595 832 676 865
rect -145 745 -111 779
rect 1384 745 1418 779
rect -146 16 -112 50
rect 1384 12 1418 46
rect 591 -38 674 -25
rect 591 -72 674 -38
rect 591 -83 674 -72
<< metal1 >>
rect 583 870 690 876
rect 583 859 595 870
rect 270 832 595 859
rect 676 859 690 870
rect 676 832 1008 859
rect 270 826 1008 832
rect -189 779 -67 785
rect -189 745 -145 779
rect -111 745 -67 779
rect -189 739 -67 745
rect -189 689 -155 739
rect -101 694 -67 739
rect -101 689 29 694
rect -84 522 29 689
rect -84 518 46 522
rect 12 474 46 518
rect 12 428 74 474
rect -121 364 -111 416
rect -59 364 -49 416
rect -102 276 -68 364
rect -85 101 28 276
rect -190 56 -156 101
rect -102 100 28 101
rect -102 56 -68 100
rect -190 50 -68 56
rect -190 16 -146 50
rect -112 16 -68 50
rect -190 10 -68 16
rect 270 -62 300 826
rect 585 706 690 826
rect 344 474 378 525
rect 344 428 406 474
rect 328 100 338 152
rect 390 100 400 152
rect 579 100 693 706
rect 872 642 882 694
rect 934 642 944 694
rect 865 320 928 366
rect 894 268 928 320
rect 579 -19 685 100
rect 579 -25 686 -19
rect 579 -29 591 -25
rect 582 -62 591 -29
rect 579 -83 591 -62
rect 674 -29 686 -25
rect 977 -28 1008 826
rect 1340 779 1462 785
rect 1340 745 1384 779
rect 1418 745 1462 779
rect 1340 739 1462 745
rect 1340 706 1374 739
rect 1428 706 1462 739
rect 1243 522 1356 694
rect 1243 518 1374 522
rect 1340 434 1374 518
rect 1321 382 1331 434
rect 1383 382 1393 434
rect 1197 320 1260 366
rect 1226 276 1260 320
rect 1226 268 1356 276
rect 1243 100 1356 268
rect 1340 52 1374 88
rect 1428 52 1462 88
rect 1340 46 1462 52
rect 1340 12 1384 46
rect 1418 12 1462 46
rect 1340 6 1462 12
rect 969 -29 1008 -28
rect 674 -62 1008 -29
rect 674 -83 686 -62
rect 579 -89 686 -83
<< rmetal1 >>
rect 300 -62 582 -29
<< via1 >>
rect -111 364 -59 416
rect 338 100 390 152
rect 882 642 934 694
rect 1331 382 1383 434
<< metal2 >>
rect 882 694 934 704
rect -111 416 -59 426
rect 339 416 391 417
rect 882 416 934 642
rect 1331 434 1383 444
rect -59 382 1331 416
rect -59 381 1383 382
rect -111 354 -59 364
rect 339 162 391 381
rect 1331 372 1383 381
rect 338 153 391 162
rect 338 152 390 153
rect 338 90 390 100
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1729327062
transform 1 0 1401 0 1 188
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1729327062
transform 1 0 -129 0 1 188
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1729327062
transform 1 0 -128 0 1 606
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1729327062
transform 1 0 1401 0 1 606
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_C77M8X  sky130_fd_pr__nfet_01v8_C77M8X_0
timestamp 1729327062
transform 1 0 636 0 1 397
box -636 -397 636 397
<< labels >>
flabel viali 623 851 623 851 0 FreeSans 1120 0 0 0 gnd
port 0 nsew
flabel metal1 26 482 26 482 0 FreeSans 1120 0 0 0 d8
port 1 nsew
flabel metal2 1279 390 1279 390 0 FreeSans 1120 0 0 0 d9
port 2 nsew
<< end >>
