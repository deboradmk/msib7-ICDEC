magic
tech sky130A
magscale 1 2
timestamp 1729427071
<< nwell >>
rect 10244 2218 11038 5118
<< metal1 >>
rect 9795 5216 9805 5225
rect 7933 5139 9805 5216
rect 7933 5054 7999 5139
rect 9795 5130 9805 5139
rect 9944 5216 9954 5225
rect 9944 5139 10608 5216
rect 9944 5130 9954 5139
rect 7933 5052 7967 5054
rect 8114 4684 8174 4690
rect 8174 4624 8428 4684
rect 8114 4618 8174 4624
rect 10527 4467 10608 5139
rect 10560 4464 10608 4467
rect 7946 4300 8138 4303
rect 7812 4267 8138 4300
rect 7812 4264 7996 4267
rect 8104 3871 8138 4267
rect 8104 3835 8335 3871
rect 8975 3768 9067 3876
rect 8981 3479 9066 3768
rect 10244 3730 10614 3778
rect 8981 3394 9225 3479
rect 10410 3451 10429 3497
rect 9118 3187 9225 3394
rect 10340 3387 10429 3451
rect 10341 3355 10429 3387
rect 9634 3317 10429 3355
rect 9634 3278 10415 3317
rect 9140 3154 9194 3187
rect 9634 3071 9711 3278
rect 10341 3250 10415 3278
<< via1 >>
rect 9805 5130 9944 5225
rect 8114 4624 8174 4684
<< metal2 >>
rect 9805 5225 9944 5235
rect 9805 5120 9944 5130
rect 8116 4684 8172 4691
rect 8108 4624 8114 4684
rect 8174 4624 8180 4684
rect 8116 4617 8172 4624
rect 9090 4398 9788 4460
rect 10928 4049 11030 4139
rect 7803 3642 7812 3702
rect 7872 3642 7881 3702
rect 8330 3672 8484 3682
rect 7334 3604 7392 3620
rect 7334 3568 7434 3604
rect 7944 3576 8330 3640
rect 7334 3122 7392 3568
rect 8330 3538 8484 3548
rect 10138 3198 10330 3208
rect 10138 3032 10330 3042
rect 9872 2796 9970 2848
rect 8375 2610 8443 2741
rect 9918 2702 9970 2796
rect 8374 2332 8443 2610
rect 9907 2394 9975 2702
rect 9892 2384 9986 2394
rect 9892 2294 9986 2304
<< via2 >>
rect 8116 4626 8172 4682
rect 7812 3642 7872 3702
rect 8330 3548 8484 3672
rect 10138 3042 10330 3198
rect 9892 2304 9986 2384
<< metal3 >>
rect 8111 4682 8177 4687
rect 8111 4626 8116 4682
rect 8172 4626 8177 4682
rect 8111 4621 8177 4626
rect 7807 3702 7877 3707
rect 8114 3702 8174 4621
rect 8505 4444 8575 4449
rect 8505 4384 8510 4444
rect 8570 4384 8575 4444
rect 8505 4379 8575 4384
rect 7807 3642 7812 3702
rect 7872 3642 8174 3702
rect 8320 3672 10129 3677
rect 7807 3637 7877 3642
rect 8320 3548 8330 3672
rect 8484 3548 10129 3672
rect 8320 3544 10129 3548
rect 8320 3543 8494 3544
rect 10000 3468 10129 3544
rect 9999 3367 10775 3468
rect 10128 3198 10340 3203
rect 10128 3042 10138 3198
rect 10330 3042 10340 3198
rect 10128 3037 10340 3042
rect 9882 2387 9996 2389
rect 9877 2384 9996 2387
rect 9877 2304 9892 2384
rect 9986 2378 9996 2384
rect 10181 2378 10285 3037
rect 9986 2304 10952 2378
rect 9877 2297 10952 2304
use nmoscs2  nmoscs2_0
timestamp 1729344768
transform 1 0 8541 0 1 2415
box -290 -89 1590 876
use nmoscs  nmoscs_0
timestamp 1729346748
transform 1 0 8622 0 1 3824
box -386 -78 1166 1266
use pmoscs2  pmoscs2_0
timestamp 1729408806
transform 1 0 10420 0 1 2522
box -176 -305 622 2014
use pmoscs  pmoscs_0
timestamp 1729246295
transform 1 0 7256 0 1 3509
box -186 -1295 868 1613
<< labels >>
flabel metal1 10025 5154 10025 5154 0 FreeSans 1120 0 0 0 vdd
port 0 nsew
flabel metal2 11019 4107 11019 4107 0 FreeSans 1120 0 0 0 vip
port 1 nsew
flabel metal2 9723 4411 9723 4411 0 FreeSans 1120 0 0 0 rs
port 2 nsew
flabel metal1 10263 3755 10263 3755 0 FreeSans 1120 0 0 0 vin
port 3 nsew
flabel metal3 10214 2354 10214 2354 0 FreeSans 1120 0 0 0 out
port 4 nsew
flabel metal1 9137 3420 9137 3420 0 FreeSans 1120 0 0 0 gnd
port 5 nsew
<< end >>
